----------------------------------------------------------------------
-- Authors: Akram Atassi and Adam Dia
-- Name: template.vhd
-- Description: template file
----------------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

entity template is
    port(
        i_in : in std_logic;
        o_out : out std_logic);
end template;

architecture rtl of template is
-- Signals

    begin


end rtl;